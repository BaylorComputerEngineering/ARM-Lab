`timescale 1ns / 1ps
`define CYCLE 10
`define WORD  64
`define INSTR_LEN 32
`define DMEMFILE  "H:/ELC3338/Spring2018/potter/ARM-Lab/testfiles/ramData.data"
`define IMEMFILE  "H:/ELC3338/Spring2018/potter/ARM-Lab/testfiles/instrData.data"
`define RMEMFILE  "H:/ELC3338/Spring2018/potter/ARM-Lab/testfiles/regData.data"
